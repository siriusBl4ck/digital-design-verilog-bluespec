always @ (input1 or input2)
    begin
        and_gate = input1 & input2;
    end